     /*
module Instruction_Memory  (PC, instruction); 

    input       [31:0]  PC;        // Input Address 

    output   [31:0]  instruction;    // Instruction at memory location Address
    
    reg [31:0] mem[0:128];


    /* Please fill in the implementation here */
     /*

	initial
	begin
		//       6    5    5    5    5       6
		//R-type op   rs   rt   rd   shamt   funt
		//I-type op   rs   rt   adress/immediate
		//J-type op        target address
		// R  lenh rd rs rt 
		// I  lenh t s immediate
		// Br lenh s t label
		mem[0] = 32'b001000_00000_00001_0000000000000101;
		mem[1] = 32'b001000_00000_00010_0000000000000111;
		mem[2] = 32'b001000_00000_00011_0000000000001100;
		mem[3] = 32'b000000_00001_00010_00100_00000_100000;
		mem[4] = 32'b000101_00100_00011_0000000000011010;
		mem[5] = 32'b101011_00000_00011_0000000000000000;
		mem[6] = 32'b100011_00000_00101_0000000000000000;
		mem[7] = 32'b000101_00101_00011_0000000000010111;
		mem[8] = 32'b000000_00010_00001_00110_00000_100010;
		mem[9] = 32'b000100_00110_00011_0000000000010101;
		mem[10]= 32'b000000_00000_00011_00111_00110_000011;
		mem[11]= 32'b000000_00111_00011_00111_00000_100100;
		mem[12]= 32'b000000_00001_00010_00001_00000_100010;
		mem[13]= 32'b000000_00001_00111_00100_00000_100110;
		mem[14]= 32'b001110_00000_00101_0000000000000010;
		mem[15]= 32'b000000_00111_00101_00010_00000_000111;
		mem[16]= 32'b101011_00101_00100_0000000000000000;
		mem[17]= 32'b100011_00101_00110_0000000000000000;
		mem[18]= 32'b101011_00101_00011_0000000000000010;
		mem[19]= 32'b100011_00101_00111_0000000000000010;
		mem[20]= 32'b000000_00101_00111_00111_00000_100101;
		mem[21]= 32'b001100_00110_00110_0000000000001101;
		mem[22]= 32'b000101_00111_00011_0000000000001000;
		mem[23]= 32'b001000_00000_00001_0000000000000101;
		mem[24]= 32'b001000_00000_00001_0000000000000101;
		mem[25]= 32'b001000_00000_00001_0000000000000101;
		mem[26]= 32'b001000_00000_00001_0000000000000101;
		
		mem[27]= 32'b001101_00000_00010_0000000000000111;//ORI $2,$0,7 		$2=7
		mem[28]= 32'b000000_00111_00000_00001_00000_100111;//NOR $1,$7,$0 	$1=-8
		mem[29]= 32'b000000_00001_00010_00000_00000_011010;//DIV $1,$2			lo=0, hi=1
		mem[30]= 32'b000000_00001_00010_00000_00000_011000;//MULT $1,$2		lo=56, hi=0
	
     /*
		0:	Inst = 10010_001_000_00101;	//ADDI $1,$0,5  	$1=5
		1:	Inst = 10010_010_000_00111;	//ADDI $2,$0,7		$2=7 	
		2:	Inst = 10010_011_000_01100;	//ADDI $3,$0,12 	$3=12
		3:	Inst = 00010_100_001_010_00;	//ADD $4,$1,$2		$4=5+7=12
		4:	Inst = 11111_011_100_11010;	//BNE $3,$4,26		if($3!=$4) PC=PC+26
		5:	Inst = 11101_011_000_00000;	//SW $3,$0,0		MEM[0]<-$3 = 12
		6:	Inst = 11100_101_000_00000;	//LW $5,$0,0		$5=12	 $5<-MEM[0] = 12
		7:	Inst = 11111_011_101_10111;	//BNE $3,$5,23		IF($3!=$5) PC=PC+23
		8:	Inst = 00011_110_010_001_00;	//SUB $6,$2,$1		$6=7-5=2
		9: 	Inst = 11110_110_011_10101;	//BEQ $6,$3,21		IF(2==12) PC=PC+12
		10:	Inst = 01000_111_100_110_00;	//SRA $7,$3,$6		$7=12>>2=3
		11:	Inst = 00100_111_111_011_00;	//AND $7,$7,$3		$7=0;
		12:	Inst = 00011_001_001_010_00;	//SUB $1,$1,$2		$1=5-7=-2
		13:	Inst = 00110_100_001_111_00;	//XOR $4,$1,$7		$4=-2
		14:	Inst = 10110_101_000_00010;	//XORI $5,$0,2		$5=2
		15:	Inst = 01001_010_101_111_00;	//SRAV $2,$5,$7		$2=2>>>0=2
		16:	Inst = 11101_100_101_00000;	//SW $4,$5,0		MEM[2]<-$4 = -2
		17:	Inst = 11100_110_101_00000;	//LW $6,$5,0		$6=Mem[2] = -2
		18:	Inst = 11101_011_101_00010;	//SW $3,$5,2		Mem[4]<-$3 = 12
		19:	Inst = 11100_111_101_00010;	//LW $7,$5,2		$7=Mem[4] = 12
		20:	Inst = 00101_111_101_111_00;	//OR $7,$5,$7		$7=14
		21:	Inst = 10100_110_110_01101;	//ANDI $6,$6,13	$6=1101&1110
		22:	Inst = 11111_111_011_01000;	//BNE $7,$3,8		if(14!=12) PC=PC+8=22+8=30

	*/    /*
	end
	assign instruction = mem[PC>>2];	
	

endmodule		*/
module Instruction_Memory  (PC, instruction); 

    input       [31:0]  PC;        // Input Address 

    output   [31:0]  instruction;    // Instruction at memory location Address
    
    reg [31:0] mem[0:1024];


	initial
	begin
		$readmemb("code.txt",mem);
	end

	assign instruction = mem[PC>>2];	
	

endmodule
